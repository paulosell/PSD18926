-- Sistema digital baseado nos Circuitos 4 e 5. O sistema deve
-- possuir quatro entradas de requisição e três saídas. Uma saída deve ser acionada sempre
-- que pelo menos uma requisição for ativada. As outras duas saídas devem identificar a
-- requisição selecionada quando alguma delas for ativada, sendo que seu valor default é "00"

library ieee;
use ieee.std_logic_1164.all;

entity one_hot_bin_system is
  port
  (
    i_REQ       : in std_logic_vector(3 downto 0);
    o_GRANT_BIT : out std_logic;
    o_GRANT_BIN : out std_logic_vector(1 downto 0)
  );
end one_hot_bin_system;

architecture arch of one_hot_bin_system is

  component one_hot_bin is
    port
    (
      i_REQ       : in std_logic_vector(3 downto 0);
      o_GRANT     : out std_logic_vector(3 downto 0);
      o_GRANT_BIN : out std_logic_vector(1 downto 0)
    );
  end component;

	-- sinal declarado apenas para instanciar o componente
  signal w_GRANT : std_logic_vector(3 downto 0);

begin
  u_1 : one_hot_bin port map
    (i_REQ => i_REQ, o_GRANT_BIN => o_GRANT_BIN, o_GRANT => w_GRANT);
  o_GRANT_BIT <= i_REQ(0) or i_REQ(1) or i_REQ(2) or i_REQ(3);
end arch;





-- Extensão do codificador de prioridades estáticas do Circuito 4
-- que apresente o identificador da requisição selecionada utilizando codificação binária de
-- dois bits. 
library ieee;
use ieee.std_logic_1164.all;


entity one_hot_bin is
  port
  (
    i_REQ       : in std_logic_vector(3 downto 0);
    o_GRANT     : out std_logic_vector(3 downto 0);
    o_GRANT_BIN : out std_logic_vector(1 downto 0)
  );
end one_hot_bin;

architecture arch of one_hot_bin is
  -- Components declaration
  component one_hot is
    port
    (
      i_REQ   : in std_logic_vector(3 downto 0);
      o_GRANT : out std_logic_vector(3 downto 0)
    );
  end component;
begin
  process (i_REQ)
  begin
    o_GRANT_BIN <= (others => '0');
    if (i_REQ(0) = '1') then
      o_GRANT_BIN <= "00";
    elsif (i_REQ(1) = '1') then
      o_GRANT_BIN <= "01";
    elsif (i_REQ(2) = '1') then
      o_GRANT_BIN <= "10";
    elsif (i_REQ(3) = '1') then
      o_GRANT_BIN <= "11";
    end if;
  end process;

  u_1 : one_hot port map
  (
    i_REQ   => i_REQ,
    o_GRANT => o_GRANT);

end arch;


---------------- definition of one hot
library ieee;
use ieee.std_logic_1164.all;

entity one_hot is
  port
  (
    i_REQ   : in std_logic_vector(3 downto 0);
    o_GRANT : out std_logic_vector(3 downto 0)
  );
end one_hot;

architecture arch of one_hot is
begin
  process (i_REQ)
  begin
    o_GRANT <= (others => '0');
    if (i_REQ(0) = '1') then
      o_GRANT(0) <= '1';
    elsif (i_REQ(1) = '1') then
      o_GRANT(1) <= '1';
    elsif (i_REQ(2) = '1') then
      o_GRANT(2) <= '1';
    elsif (i_REQ(3) = '1') then
      o_GRANT(3) <= '1';
    end if;
  end process;
end arch;